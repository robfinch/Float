// ============================================================================
//        __
//   \\__/ o\    (C) 2020-2022  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//	mult64x64_tb.sv
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// ============================================================================

module mult64x64_tb();
reg clk;
reg [23:0] count;
reg [31:0] adr;

reg rst;
reg [63:0] a, b;
wire [127:0] o;
wire [127:0] p = a * b;

always #5 clk = ~clk;

mult64x64 u1 (clk, 1'b1, a, b, o);

integer outfile;

initial begin
	rst = 1'b0;
	clk = 1'b0;
	#20 rst = 1;
	#50 rst = 0;
	#1000000  $fclose(outfile);
	#10 $finish;
end

always #5
	clk = ~clk;

always_ff @(posedge clk)
if (rst) begin
	adr <= 0;
	count <= 0;
	a <= $urandom(1);
end
else
begin
  if (adr==0) begin
    outfile = $fopen("d:/cores2022/rf6809/rtl/fpu/test_bench/mult64x64_tvo.txt", "wb");
    $fwrite(outfile, "--- A ---  ---- B ----  - DUT Product -  - SIM Product -\n");
  end
	count <= count + 1;
	if (count > 24)
		count <= 1'd1;
	if (count==2) begin	
		case (adr)
	  1:
	    begin
	      a <= 64'd10;
	      b <= 64'd10;
	    end
	  2:
	    begin
	      a <= 64'd21;
	      b <= 64'd1700000;
	    end 
	  3:
	    begin
	      a <= 64'd215000;
	      b <= 64'd11;
	    end
	  default:
	  	begin
				a[31:0] <= $urandom();
				b[31:0] <= $urandom();
				a[63:32] <= $urandom();
				b[63:32] <= $urandom();
			end
	  endcase 
	end
	if (count==24) begin
	  $fwrite(outfile, "%h\t%h\t%h\t%h%c\n", a, b, o, p,p!=o ? "*":" ");
		adr <= adr + 1;
	end
end

endmodule
