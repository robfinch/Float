module FP2DFP128a();



endmodule

module ShiftReg(clk, adr, i, o);
input [15:0] adr;

reg [63:0] mem [0:1023];


endmodule
