// ============================================================================
//        __
//   \\__/ o\    (C) 2020-2022  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//	DFPRes128.sv
//  - estimate the reciprocal of number between 0.1 and 1.0
//  - the reciprocal is between 1.00 and 9.99
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//                                                                          
// ============================================================================

import DFPPkg::*;

module DFPRes128(clk, i, o);
input clk;
input [127:0] i;
output [127:0] o;

DFP128U iu, ou;
DFPUnpack128 u1 (i, iu);

reg [11:0] ndx;
(* ram_style = "block" *)
reg [23:0] mem [0:4095];

initial begin
	mem[16'h000] = 24'hFFFFFF; //xxxxxxxxx
	mem[16'h001] = 24'h000000; //005f5e100
	mem[16'h002] = 24'h000000; //002faf080
	mem[16'h003] = 24'h333333; //001fca055
	mem[16'h004] = 24'h000000; //0017d7840
	mem[16'h005] = 24'h000000; //001312d00
	mem[16'h006] = 24'h666666; //000fe502a
	mem[16'h007] = 24'h285714; //000d9fb92
	mem[16'h008] = 24'h500000; //000bebc20
	mem[16'h009] = 24'h111111; //000a98ac7
	mem[16'h080] = 24'h250000; //0001312d0
	mem[16'h081] = 24'h234567; //00012d687
	mem[16'h800] = 24'h125000; //00001e848
	mem[16'h801] = 24'h124843; //00001e7ab
	mem[16'h880] = 24'h113636; //00001bbe4
	mem[16'h881] = 24'h113507; //00001bb63
	mem[16'h010] = 24'h000000; //000989680
	mem[16'h011] = 24'h090909; //0008ab75d
	mem[16'h012] = 24'h333333; //0007f2815
	mem[16'h013] = 24'h692307; //000756013
	mem[16'h014] = 24'h142857; //0006cfdc9
	mem[16'h015] = 24'h666666; //00065b9aa
	mem[16'h016] = 24'h250000; //0005f5e10
	mem[16'h017] = 24'h882352; //00059c1f0
	mem[16'h018] = 24'h555555; //00054c563
	mem[16'h019] = 24'h263157; //000504f35
	mem[16'h090] = 24'h111111; //00010f447
	mem[16'h091] = 24'h098901; //00010c495
	mem[16'h810] = 24'h123456; //00001e240
	mem[16'h811] = 24'h123304; //00001e1a8
	mem[16'h890] = 24'h112359; //00001b6e7
	mem[16'h891] = 24'h112233; //00001b669
	mem[16'h020] = 24'h000000; //0004c4b40
	mem[16'h021] = 24'h761904; //00048a930
	mem[16'h022] = 24'h545454; //000455bae
	mem[16'h023] = 24'h347826; //0004257b2
	mem[16'h024] = 24'h166666; //0003f940a
	mem[16'h025] = 24'h000000; //0003d0900
	mem[16'h026] = 24'h846153; //0003ab009
	mem[16'h027] = 24'h703703; //000388397
	mem[16'h028] = 24'h571428; //000367ee4
	mem[16'h029] = 24'h448275; //000349dd3
	mem[16'h082] = 24'h219512; //000129bb8
	mem[16'h083] = 24'h204819; //000126253
	mem[16'h820] = 24'h121951; //00001dc5f
	mem[16'h821] = 24'h121802; //00001dbca
	mem[16'h808] = 24'h123762; //00001e372
	mem[16'h809] = 24'h123609; //00001e2d9
	mem[16'h030] = 24'h333333; //00032dcd5
	mem[16'h031] = 24'h225806; //0003138ce
	mem[16'h032] = 24'h125000; //0002faf08
	mem[16'h033] = 24'h030303; //0002e3d1f
	mem[16'h034] = 24'h941176; //0002ce0f8
	mem[16'h035] = 24'h857142; //0002b98b6
	mem[16'h036] = 24'h777777; //0002a62b1
	mem[16'h037] = 24'h702702; //000293d6e
	mem[16'h038] = 24'h631578; //00028279a
	mem[16'h039] = 24'h564102; //000272006
	mem[16'h092] = 24'h086956; //0001095ec
	mem[16'h093] = 24'h075268; //000106844
	mem[16'h830] = 24'h120481; //00001d6a1
	mem[16'h831] = 24'h120336; //00001d610
	mem[16'h818] = 24'h122249; //00001dd89
	mem[16'h819] = 24'h122100; //00001dcf4
	mem[16'h040] = 24'h500000; //0002625a0
	mem[16'h041] = 24'h439024; //000253770
	mem[16'h042] = 24'h380952; //000245498
	mem[16'h043] = 24'h325581; //000237c4d
	mem[16'h044] = 24'h272727; //00022add7
	mem[16'h045] = 24'h222222; //00021e88e
	mem[16'h046] = 24'h173913; //000212bd9
	mem[16'h047] = 24'h127659; //00020772b
	mem[16'h048] = 24'h083333; //0001fca05
	mem[16'h049] = 24'h040816; //0001f23f0
	mem[16'h084] = 24'h190476; //000122a4c
	mem[16'h085] = 24'h176470; //00011f396
	mem[16'h840] = 24'h119047; //00001d107
	mem[16'h841] = 24'h118906; //00001d07a
	mem[16'h088] = 24'h136363; //0001156eb
	mem[16'h089] = 24'h123595; //00011250b
	mem[16'h050] = 24'h000000; //0001e8480
	mem[16'h051] = 24'h960784; //0001deb50
	mem[16'h052] = 24'h923076; //0001d5804
	mem[16'h053] = 24'h886792; //0001cca48
	mem[16'h054] = 24'h851851; //0001c41cb
	mem[16'h055] = 24'h818181; //0001bbe45
	mem[16'h056] = 24'h785714; //0001b3f72
	mem[16'h057] = 24'h754385; //0001ac511
	mem[16'h058] = 24'h724137; //0001a4ee9
	mem[16'h059] = 24'h694915; //00019dcc3
	mem[16'h094] = 24'h063829; //000103b95
	mem[16'h095] = 24'h052631; //000100fd7
	mem[16'h850] = 24'h117647; //00001cb8f
	mem[16'h851] = 24'h117508; //00001cb04
	mem[16'h098] = 24'h020408; //0000f91f8
	mem[16'h099] = 24'h010101; //0000f69b5
	mem[16'h060] = 24'h666666; //000196e6a
	mem[16'h061] = 24'h639344; //0001903b0
	mem[16'h062] = 24'h612903; //000189c67
	mem[16'h063] = 24'h587301; //000183865
	mem[16'h064] = 24'h562500; //00017d784
	mem[16'h065] = 24'h538461; //00017799d
	mem[16'h066] = 24'h515151; //000171e8f
	mem[16'h067] = 24'h492537; //00016c639
	mem[16'h068] = 24'h470588; //00016707c
	mem[16'h069] = 24'h449275; //000161d3b
	mem[16'h086] = 24'h162790; //00011be26
	mem[16'h087] = 24'h149425; //0001189f1
	mem[16'h860] = 24'h116279; //00001c637
	mem[16'h861] = 24'h116144; //00001c5b0
	mem[16'h888] = 24'h112612; //00001b7e4
	mem[16'h889] = 24'h112485; //00001b765
	mem[16'h070] = 24'h428571; //00015cc5b
	mem[16'h071] = 24'h408450; //000157dc2
	mem[16'h072] = 24'h388888; //000153158
	mem[16'h073] = 24'h369863; //00014e707
	mem[16'h074] = 24'h351351; //000149eb7
	mem[16'h075] = 24'h333333; //000145855
	mem[16'h076] = 24'h315789; //0001413cd
	mem[16'h077] = 24'h298701; //00013d10d
	mem[16'h078] = 24'h282051; //000139003
	mem[16'h079] = 24'h265822; //00013509e
	mem[16'h096] = 24'h041666; //0000fe502
	mem[16'h097] = 24'h030927; //0000fbb0f
	mem[16'h870] = 24'h114942; //00001c0fe
	mem[16'h871] = 24'h114810; //00001c07a
	mem[16'h898] = 24'h111358; //00001b2fe
	mem[16'h899] = 24'h111234; //00001b282
	mem[16'h100] = 24'h999999; //0000f4240
	mem[16'h101] = 24'h990099; //0000f1b93
	mem[16'h102] = 24'h980392; //0000ef5a8
	mem[16'h103] = 24'h970873; //0000ed079
	mem[16'h104] = 24'h961538; //0000eac02
	mem[16'h105] = 24'h952380; //0000e883c
	mem[16'h106] = 24'h943396; //0000e6524
	mem[16'h107] = 24'h934579; //0000e42b3
	mem[16'h108] = 24'h925925; //0000e20e5
	mem[16'h109] = 24'h917431; //0000dffb7
	mem[16'h180] = 24'h555555; //000087a23
	mem[16'h181] = 24'h552486; //000086e26
	mem[16'h900] = 24'h111111; //00001b207
	mem[16'h901] = 24'h110987; //00001b18b
	mem[16'h980] = 24'h102040; //000018e98
	mem[16'h981] = 24'h101936; //000018e30
	mem[16'h110] = 24'h909090; //0000ddf22
	mem[16'h111] = 24'h900900; //0000dbf24
	mem[16'h112] = 24'h892857; //0000d9fb9
	mem[16'h113] = 24'h884955; //0000d80db
	mem[16'h114] = 24'h877192; //0000d6288
	mem[16'h115] = 24'h869565; //0000d44bd
	mem[16'h116] = 24'h862068; //0000d2774
	mem[16'h117] = 24'h854700; //0000d0aac
	mem[16'h118] = 24'h847457; //0000cee61
	mem[16'h119] = 24'h840336; //0000cd290
	mem[16'h190] = 24'h526315; //0000807eb
	mem[16'h191] = 24'h523560; //00007fd28
	mem[16'h910] = 24'h109890; //00001ad42
	mem[16'h911] = 24'h109769; //00001acc9
	mem[16'h990] = 24'h101010; //000018a92
	mem[16'h991] = 24'h100908; //000018a2c
	mem[16'h120] = 24'h833333; //0000cb735
	mem[16'h121] = 24'h826446; //0000c9c4e
	mem[16'h122] = 24'h819672; //0000c81d8
	mem[16'h123] = 24'h813008; //0000c67d0
	mem[16'h124] = 24'h806451; //0000c4e33
	mem[16'h125] = 24'h800000; //0000c3500
	mem[16'h126] = 24'h793650; //0000c1c32
	mem[16'h127] = 24'h787401; //0000c03c9
	mem[16'h128] = 24'h781250; //0000bebc2
	mem[16'h129] = 24'h775193; //0000bd419
	mem[16'h182] = 24'h549450; //00008624a
	mem[16'h183] = 24'h546448; //000085690
	mem[16'h920] = 24'h108695; //00001a897
	mem[16'h921] = 24'h108577; //00001a821
	mem[16'h908] = 24'h110132; //00001ae34
	mem[16'h909] = 24'h110011; //00001adbb
	mem[16'h130] = 24'h769230; //0000bbcce
	mem[16'h131] = 24'h763358; //0000ba5de
	mem[16'h132] = 24'h757575; //0000b8f47
	mem[16'h133] = 24'h751879; //0000b7907
	mem[16'h134] = 24'h746268; //0000b631c
	mem[16'h135] = 24'h740740; //0000b4d84
	mem[16'h136] = 24'h735294; //0000b383e
	mem[16'h137] = 24'h729927; //0000b2347
	mem[16'h138] = 24'h724637; //0000b0e9d
	mem[16'h139] = 24'h719424; //0000afa40
	mem[16'h192] = 24'h520833; //00007f281
	mem[16'h193] = 24'h518134; //00007e7f6
	mem[16'h930] = 24'h107526; //00001a406
	mem[16'h931] = 24'h107411; //00001a393
	mem[16'h918] = 24'h108932; //00001a984
	mem[16'h919] = 24'h108813; //00001a90d
	mem[16'h140] = 24'h714285; //0000ae62d
	mem[16'h141] = 24'h709219; //0000ad263
	mem[16'h142] = 24'h704225; //0000abee1
	mem[16'h143] = 24'h699300; //0000aaba4
	mem[16'h144] = 24'h694444; //0000a98ac
	mem[16'h145] = 24'h689655; //0000a85f7
	mem[16'h146] = 24'h684931; //0000a7383
	mem[16'h147] = 24'h680272; //0000a6150
	mem[16'h148] = 24'h675675; //0000a4f5b
	mem[16'h149] = 24'h671140; //0000a3da4
	mem[16'h184] = 24'h543478; //000084af6
	mem[16'h185] = 24'h540540; //000083f7c
	mem[16'h940] = 24'h106382; //000019f8e
	mem[16'h941] = 24'h106269; //000019f1d
	mem[16'h188] = 24'h531914; //000081dca
	mem[16'h189] = 24'h529100; //0000812cc
	mem[16'h150] = 24'h666666; //0000a2c2a
	mem[16'h151] = 24'h662251; //0000a1aeb
	mem[16'h152] = 24'h657894; //0000a09e6
	mem[16'h153] = 24'h653594; //00009f91a
	mem[16'h154] = 24'h649350; //00009e886
	mem[16'h155] = 24'h645161; //00009d829
	mem[16'h156] = 24'h641025; //00009c801
	mem[16'h157] = 24'h636942; //00009b80e
	mem[16'h158] = 24'h632911; //00009a84f
	mem[16'h159] = 24'h628930; //0000998c2
	mem[16'h194] = 24'h515463; //00007dd87
	mem[16'h195] = 24'h512820; //00007d334
	mem[16'h950] = 24'h105263; //000019b2f
	mem[16'h951] = 24'h105152; //000019ac0
	mem[16'h198] = 24'h505050; //00007b4da
	mem[16'h199] = 24'h502512; //00007aaf0
	mem[16'h160] = 24'h625000; //000098968
	mem[16'h161] = 24'h621118; //000097a3e
	mem[16'h162] = 24'h617283; //000096b43
	mem[16'h163] = 24'h613496; //000095c78
	mem[16'h164] = 24'h609756; //000094ddc
	mem[16'h165] = 24'h606060; //000093f6c
	mem[16'h166] = 24'h602409; //000093129
	mem[16'h167] = 24'h598802; //000092312
	mem[16'h168] = 24'h595238; //000091526
	mem[16'h169] = 24'h591715; //000090763
	mem[16'h186] = 24'h537634; //000083422
	mem[16'h187] = 24'h534759; //0000828e7
	mem[16'h960] = 24'h104166; //0000196e6
	mem[16'h961] = 24'h104058; //00001967a
	mem[16'h988] = 24'h101214; //000018b5e
	mem[16'h989] = 24'h101112; //000018af8
	mem[16'h170] = 24'h588235; //00008f9cb
	mem[16'h171] = 24'h584795; //00008ec5b
	mem[16'h172] = 24'h581395; //00008df13
	mem[16'h173] = 24'h578034; //00008d1f2
	mem[16'h174] = 24'h574712; //00008c4f8
	mem[16'h175] = 24'h571428; //00008b824
	mem[16'h176] = 24'h568181; //00008ab75
	mem[16'h177] = 24'h564971; //000089eeb
	mem[16'h178] = 24'h561797; //000089285
	mem[16'h179] = 24'h558659; //000088643
	mem[16'h196] = 24'h510204; //00007c8fc
	mem[16'h197] = 24'h507614; //00007bede
	mem[16'h970] = 24'h103092; //0000192b4
	mem[16'h971] = 24'h102986; //00001924a
	mem[16'h998] = 24'h100200; //000018768
	mem[16'h999] = 24'h100100; //000018704
	mem[16'h200] = 24'h500000; //00007a120
	mem[16'h201] = 24'h497512; //000079768
	mem[16'h202] = 24'h495049; //000078dc9
	mem[16'h203] = 24'h492610; //000078442
	mem[16'h204] = 24'h490196; //000077ad4
	mem[16'h205] = 24'h487804; //00007717c
	mem[16'h206] = 24'h485436; //00007683c
	mem[16'h207] = 24'h483091; //000075f13
	mem[16'h208] = 24'h480769; //000075601
	mem[16'h209] = 24'h478468; //000074d04
	mem[16'h280] = 24'h357142; //000057316
	mem[16'h281] = 24'h355871; //000056e1f
	mem[16'h802] = 24'h124688; //00001e710
	mem[16'h803] = 24'h124533; //00001e675
	mem[16'h882] = 24'h113378; //00001bae2
	mem[16'h883] = 24'h113250; //00001ba62
	mem[16'h210] = 24'h476190; //00007441e
	mem[16'h211] = 24'h473933; //000073b4d
	mem[16'h212] = 24'h471698; //000073292
	mem[16'h213] = 24'h469483; //0000729eb
	mem[16'h214] = 24'h467289; //000072159
	mem[16'h215] = 24'h465116; //0000718dc
	mem[16'h216] = 24'h462962; //000071072
	mem[16'h217] = 24'h460829; //00007081d
	mem[16'h218] = 24'h458715; //00006ffdb
	mem[16'h219] = 24'h456621; //00006f7ad
	mem[16'h290] = 24'h344827; //0000542fb
	mem[16'h291] = 24'h343642; //000053e5a
	mem[16'h812] = 24'h123152; //00001e110
	mem[16'h813] = 24'h123001; //00001e079
	mem[16'h892] = 24'h112107; //00001b5eb
	mem[16'h893] = 24'h111982; //00001b56e
	mem[16'h220] = 24'h454545; //00006ef91
	mem[16'h221] = 24'h452488; //00006e788
	mem[16'h222] = 24'h450450; //00006df92
	mem[16'h223] = 24'h448430; //00006d7ae
	mem[16'h224] = 24'h446428; //00006cfdc
	mem[16'h225] = 24'h444444; //00006c81c
	mem[16'h226] = 24'h442477; //00006c06d
	mem[16'h227] = 24'h440528; //00006b8d0
	mem[16'h228] = 24'h438596; //00006b144
	mem[16'h229] = 24'h436681; //00006a9c9
	mem[16'h282] = 24'h354609; //000056931
	mem[16'h283] = 24'h353356; //00005644c
	mem[16'h822] = 24'h121654; //00001db36
	mem[16'h823] = 24'h121506; //00001daa2
	mem[16'h828] = 24'h120772; //00001d7c4
	mem[16'h829] = 24'h120627; //00001d733
	mem[16'h230] = 24'h434782; //00006a25e
	mem[16'h231] = 24'h432900; //000069b04
	mem[16'h232] = 24'h431034; //0000693ba
	mem[16'h233] = 24'h429184; //000068c80
	mem[16'h234] = 24'h427350; //000068556
	mem[16'h235] = 24'h425531; //000067e3b
	mem[16'h236] = 24'h423728; //000067730
	mem[16'h237] = 24'h421940; //000067034
	mem[16'h238] = 24'h420168; //000066948
	mem[16'h239] = 24'h418410; //00006626a
	mem[16'h292] = 24'h342465; //0000539c1
	mem[16'h293] = 24'h341296; //000053530
	mem[16'h832] = 24'h120192; //00001d580
	mem[16'h833] = 24'h120048; //00001d4f0
	mem[16'h838] = 24'h119331; //00001d223
	mem[16'h839] = 24'h119189; //00001d195
	mem[16'h240] = 24'h416666; //000065b9a
	mem[16'h241] = 24'h414937; //0000654d9
	mem[16'h242] = 24'h413223; //000064e27
	mem[16'h243] = 24'h411522; //000064782
	mem[16'h244] = 24'h409836; //0000640ec
	mem[16'h245] = 24'h408163; //000063a63
	mem[16'h246] = 24'h406504; //0000633e8
	mem[16'h247] = 24'h404858; //000062d7a
	mem[16'h248] = 24'h403225; //000062719
	mem[16'h249] = 24'h401606; //0000620c6
	mem[16'h284] = 24'h352112; //000055f70
	mem[16'h285] = 24'h350877; //000055a9d
	mem[16'h842] = 24'h118764; //00001cfec
	mem[16'h843] = 24'h118623; //00001cf5f
	mem[16'h288] = 24'h347222; //000054c56
	mem[16'h289] = 24'h346020; //0000547a4
	mem[16'h250] = 24'h400000; //000061a80
	mem[16'h251] = 24'h398406; //000061446
	mem[16'h252] = 24'h396825; //000060e19
	mem[16'h253] = 24'h395256; //0000607f8
	mem[16'h254] = 24'h393700; //0000601e4
	mem[16'h255] = 24'h392156; //00005fbdc
	mem[16'h256] = 24'h390625; //00005f5e1
	mem[16'h257] = 24'h389105; //00005eff1
	mem[16'h258] = 24'h387596; //00005ea0c
	mem[16'h259] = 24'h386100; //00005e434
	mem[16'h294] = 24'h340136; //0000530a8
	mem[16'h295] = 24'h338983; //000052c27
	mem[16'h852] = 24'h117370; //00001ca7a
	mem[16'h853] = 24'h117233; //00001c9f1
	mem[16'h298] = 24'h335570; //000051ed2
	mem[16'h299] = 24'h334448; //000051a70
	mem[16'h260] = 24'h384615; //00005de67
	mem[16'h261] = 24'h383141; //00005d8a5
	mem[16'h262] = 24'h381679; //00005d2ef
	mem[16'h263] = 24'h380228; //00005cd44
	mem[16'h264] = 24'h378787; //00005c7a3
	mem[16'h265] = 24'h377358; //00005c20e
	mem[16'h266] = 24'h375939; //00005bc83
	mem[16'h267] = 24'h374531; //00005b703
	mem[16'h268] = 24'h373134; //00005b18e
	mem[16'h269] = 24'h371747; //00005ac23
	mem[16'h286] = 24'h349650; //0000555d2
	mem[16'h287] = 24'h348432; //000055110
	mem[16'h862] = 24'h116009; //00001c529
	mem[16'h863] = 24'h115874; //00001c4a2
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h270] = 24'h370370; //00005a6c2
	mem[16'h271] = 24'h369003; //00005a16b
	mem[16'h272] = 24'h367647; //000059c1f
	mem[16'h273] = 24'h366300; //0000596dc
	mem[16'h274] = 24'h364963; //0000591a3
	mem[16'h275] = 24'h363636; //000058c74
	mem[16'h276] = 24'h362318; //00005874e
	mem[16'h277] = 24'h361010; //000058232
	mem[16'h278] = 24'h359712; //000057d20
	mem[16'h279] = 24'h358422; //000057816
	mem[16'h296] = 24'h337837; //0000527ad
	mem[16'h297] = 24'h336700; //00005233c
	mem[16'h872] = 24'h114678; //00001bff6
	mem[16'h873] = 24'h114547; //00001bf73
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h300] = 24'h333333; //000051615
	mem[16'h301] = 24'h332225; //0000511c1
	mem[16'h302] = 24'h331125; //000050d75
	mem[16'h303] = 24'h330033; //000050931
	mem[16'h304] = 24'h328947; //0000504f3
	mem[16'h305] = 24'h327868; //0000500bc
	mem[16'h306] = 24'h326797; //00004fc8d
	mem[16'h307] = 24'h325732; //00004f864
	mem[16'h308] = 24'h324675; //00004f443
	mem[16'h309] = 24'h323624; //00004f028
	mem[16'h380] = 24'h263157; //0000403f5
	mem[16'h381] = 24'h262467; //000040143
	mem[16'h902] = 24'h110864; //00001b110
	mem[16'h903] = 24'h110741; //00001b095
	mem[16'h982] = 24'h101832; //000018dc8
	mem[16'h983] = 24'h101729; //000018d61
	mem[16'h310] = 24'h322580; //00004ec14
	mem[16'h311] = 24'h321543; //00004e807
	mem[16'h312] = 24'h320512; //00004e400
	mem[16'h313] = 24'h319488; //00004e000
	mem[16'h314] = 24'h318471; //00004dc07
	mem[16'h315] = 24'h317460; //00004d814
	mem[16'h316] = 24'h316455; //00004d427
	mem[16'h317] = 24'h315457; //00004d041
	mem[16'h318] = 24'h314465; //00004cc61
	mem[16'h319] = 24'h313479; //00004c887
	mem[16'h390] = 24'h256410; //00003e99a
	mem[16'h391] = 24'h255754; //00003e70a
	mem[16'h912] = 24'h109649; //00001ac51
	mem[16'h913] = 24'h109529; //00001abd9
	mem[16'h992] = 24'h100806; //0000189c6
	mem[16'h993] = 24'h100704; //000018960
	mem[16'h320] = 24'h312500; //00004c4b4
	mem[16'h321] = 24'h311526; //00004c0e6
	mem[16'h322] = 24'h310559; //00004bd1f
	mem[16'h323] = 24'h309597; //00004b95d
	mem[16'h324] = 24'h308641; //00004b5a1
	mem[16'h325] = 24'h307692; //00004b1ec
	mem[16'h326] = 24'h306748; //00004ae3c
	mem[16'h327] = 24'h305810; //00004aa92
	mem[16'h328] = 24'h304878; //00004a6ee
	mem[16'h329] = 24'h303951; //00004a34f
	mem[16'h382] = 24'h261780; //00003fe94
	mem[16'h383] = 24'h261096; //00003fbe8
	mem[16'h922] = 24'h108459; //00001a7ab
	mem[16'h923] = 24'h108342; //00001a736
	mem[16'h928] = 24'h107758; //00001a4ee
	mem[16'h929] = 24'h107642; //00001a47a
	mem[16'h330] = 24'h303030; //000049fb6
	mem[16'h331] = 24'h302114; //000049c22
	mem[16'h332] = 24'h301204; //000049894
	mem[16'h333] = 24'h300300; //00004950c
	mem[16'h334] = 24'h299401; //000049189
	mem[16'h335] = 24'h298507; //000048e0b
	mem[16'h336] = 24'h297619; //000048a93
	mem[16'h337] = 24'h296735; //00004871f
	mem[16'h338] = 24'h295857; //0000483b1
	mem[16'h339] = 24'h294985; //000048049
	mem[16'h392] = 24'h255102; //00003e47e
	mem[16'h393] = 24'h254452; //00003e1f4
	mem[16'h932] = 24'h107296; //00001a320
	mem[16'h933] = 24'h107181; //00001a2ad
	mem[16'h938] = 24'h106609; //00001a071
	mem[16'h939] = 24'h106496; //00001a000
	mem[16'h340] = 24'h294117; //000047ce5
	mem[16'h341] = 24'h293255; //000047987
	mem[16'h342] = 24'h292397; //00004762d
	mem[16'h343] = 24'h291545; //0000472d9
	mem[16'h344] = 24'h290697; //000046f89
	mem[16'h345] = 24'h289855; //000046c3f
	mem[16'h346] = 24'h289017; //0000468f9
	mem[16'h347] = 24'h288184; //0000465b8
	mem[16'h348] = 24'h287356; //00004627c
	mem[16'h349] = 24'h286532; //000045f44
	mem[16'h384] = 24'h260416; //00003f940
	mem[16'h385] = 24'h259740; //00003f69c
	mem[16'h942] = 24'h106157; //000019ead
	mem[16'h943] = 24'h106044; //000019e3c
	mem[16'h388] = 24'h257731; //00003eec3
	mem[16'h389] = 24'h257069; //00003ec2d
	mem[16'h350] = 24'h285714; //000045c12
	mem[16'h351] = 24'h284900; //0000458e4
	mem[16'h352] = 24'h284090; //0000455ba
	mem[16'h353] = 24'h283286; //000045296
	mem[16'h354] = 24'h282485; //000044f75
	mem[16'h355] = 24'h281690; //000044c5a
	mem[16'h356] = 24'h280898; //000044942
	mem[16'h357] = 24'h280112; //000044630
	mem[16'h358] = 24'h279329; //000044321
	mem[16'h359] = 24'h278551; //000044017
	mem[16'h394] = 24'h253807; //00003df6f
	mem[16'h395] = 24'h253164; //00003dcec
	mem[16'h952] = 24'h105042; //000019a52
	mem[16'h953] = 24'h104931; //0000199e3
	mem[16'h398] = 24'h251256; //00003d578
	mem[16'h399] = 24'h250626; //00003d302
	mem[16'h360] = 24'h277777; //000043d11
	mem[16'h361] = 24'h277008; //000043a10
	mem[16'h362] = 24'h276243; //000043713
	mem[16'h363] = 24'h275482; //00004341a
	mem[16'h364] = 24'h274725; //000043125
	mem[16'h365] = 24'h273972; //000042e34
	mem[16'h366] = 24'h273224; //000042b48
	mem[16'h367] = 24'h272479; //00004285f
	mem[16'h368] = 24'h271739; //00004257b
	mem[16'h369] = 24'h271002; //00004229a
	mem[16'h386] = 24'h259067; //00003f3fb
	mem[16'h387] = 24'h258397; //00003f15d
	mem[16'h962] = 24'h103950; //00001960e
	mem[16'h963] = 24'h103842; //0000195a2
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h370] = 24'h270270; //000041fbe
	mem[16'h371] = 24'h269541; //000041ce5
	mem[16'h372] = 24'h268817; //000041a11
	mem[16'h373] = 24'h268096; //000041740
	mem[16'h374] = 24'h267379; //000041473
	mem[16'h375] = 24'h266666; //0000411aa
	mem[16'h376] = 24'h265957; //000040ee5
	mem[16'h377] = 24'h265251; //000040c23
	mem[16'h378] = 24'h264550; //000040966
	mem[16'h379] = 24'h263852; //0000406ac
	mem[16'h396] = 24'h252525; //00003da6d
	mem[16'h397] = 24'h251889; //00003d7f1
	mem[16'h972] = 24'h102880; //0000191e0
	mem[16'h973] = 24'h102774; //000019176
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h400] = 24'h250000; //00003d090
	mem[16'h401] = 24'h249376; //00003ce20
	mem[16'h402] = 24'h248756; //00003cbb4
	mem[16'h403] = 24'h248138; //00003c94a
	mem[16'h404] = 24'h247524; //00003c6e4
	mem[16'h405] = 24'h246913; //00003c481
	mem[16'h406] = 24'h246305; //00003c221
	mem[16'h407] = 24'h245700; //00003bfc4
	mem[16'h408] = 24'h245098; //00003bd6a
	mem[16'h409] = 24'h244498; //00003bb12
	mem[16'h480] = 24'h208333; //000032dcd
	mem[16'h481] = 24'h207900; //000032c1c
	mem[16'h804] = 24'h124378; //00001e5da
	mem[16'h805] = 24'h124223; //00001e53f
	mem[16'h884] = 24'h113122; //00001b9e2
	mem[16'h885] = 24'h112994; //00001b962
	mem[16'h410] = 24'h243902; //00003b8be
	mem[16'h411] = 24'h243309; //00003b66d
	mem[16'h412] = 24'h242718; //00003b41e
	mem[16'h413] = 24'h242130; //00003b1d2
	mem[16'h414] = 24'h241545; //00003af89
	mem[16'h415] = 24'h240963; //00003ad43
	mem[16'h416] = 24'h240384; //00003ab00
	mem[16'h417] = 24'h239808; //00003a8c0
	mem[16'h418] = 24'h239234; //00003a682
	mem[16'h419] = 24'h238663; //00003a447
	mem[16'h490] = 24'h204081; //000031d31
	mem[16'h491] = 24'h203665; //000031b91
	mem[16'h814] = 24'h122850; //00001dfe2
	mem[16'h815] = 24'h122699; //00001df4b
	mem[16'h894] = 24'h111856; //00001b4f0
	mem[16'h895] = 24'h111731; //00001b473
	mem[16'h420] = 24'h238095; //00003a20f
	mem[16'h421] = 24'h237529; //000039fd9
	mem[16'h422] = 24'h236966; //000039da6
	mem[16'h423] = 24'h236406; //000039b76
	mem[16'h424] = 24'h235849; //000039949
	mem[16'h425] = 24'h235294; //00003971e
	mem[16'h426] = 24'h234741; //0000394f5
	mem[16'h427] = 24'h234192; //0000392d0
	mem[16'h428] = 24'h233644; //0000390ac
	mem[16'h429] = 24'h233100; //000038e8c
	mem[16'h482] = 24'h207468; //000032a6c
	mem[16'h483] = 24'h207039; //0000328bf
	mem[16'h824] = 24'h121359; //00001da0f
	mem[16'h825] = 24'h121212; //00001d97c
	mem[16'h848] = 24'h117924; //00001cca4
	mem[16'h849] = 24'h117785; //00001cc19
	mem[16'h430] = 24'h232558; //000038c6e
	mem[16'h431] = 24'h232018; //000038a52
	mem[16'h432] = 24'h231481; //000038839
	mem[16'h433] = 24'h230946; //000038622
	mem[16'h434] = 24'h230414; //00003840e
	mem[16'h435] = 24'h229885; //0000381fd
	mem[16'h436] = 24'h229357; //000037fed
	mem[16'h437] = 24'h228832; //000037de0
	mem[16'h438] = 24'h228310; //000037bd6
	mem[16'h439] = 24'h227790; //0000379ce
	mem[16'h492] = 24'h203252; //0000319f4
	mem[16'h493] = 24'h202839; //000031857
	mem[16'h834] = 24'h119904; //00001d460
	mem[16'h835] = 24'h119760; //00001d3d0
	mem[16'h858] = 24'h116550; //00001c746
	mem[16'h859] = 24'h116414; //00001c6be
	mem[16'h440] = 24'h227272; //0000377c8
	mem[16'h441] = 24'h226757; //0000375c5
	mem[16'h442] = 24'h226244; //0000373c4
	mem[16'h443] = 24'h225733; //0000371c5
	mem[16'h444] = 24'h225225; //000036fc9
	mem[16'h445] = 24'h224719; //000036dcf
	mem[16'h446] = 24'h224215; //000036bd7
	mem[16'h447] = 24'h223713; //0000369e1
	mem[16'h448] = 24'h223214; //0000367ee
	mem[16'h449] = 24'h222717; //0000365fd
	mem[16'h484] = 24'h206611; //000032713
	mem[16'h485] = 24'h206185; //000032569
	mem[16'h844] = 24'h118483; //00001ced3
	mem[16'h845] = 24'h118343; //00001ce47
	mem[16'h488] = 24'h204918; //000032076
	mem[16'h489] = 24'h204498; //000031ed2
	mem[16'h450] = 24'h222222; //00003640e
	mem[16'h451] = 24'h221729; //000036221
	mem[16'h452] = 24'h221238; //000036036
	mem[16'h453] = 24'h220750; //000035e4e
	mem[16'h454] = 24'h220264; //000035c68
	mem[16'h455] = 24'h219780; //000035a84
	mem[16'h456] = 24'h219298; //0000358a2
	mem[16'h457] = 24'h218818; //0000356c2
	mem[16'h458] = 24'h218340; //0000354e4
	mem[16'h459] = 24'h217864; //000035308
	mem[16'h494] = 24'h202429; //0000316bd
	mem[16'h495] = 24'h202020; //000031524
	mem[16'h854] = 24'h117096; //00001c968
	mem[16'h855] = 24'h116959; //00001c8df
	mem[16'h498] = 24'h200803; //000031063
	mem[16'h499] = 24'h200400; //000030ed0
	mem[16'h460] = 24'h217391; //00003512f
	mem[16'h461] = 24'h216919; //000034f57
	mem[16'h462] = 24'h216450; //000034d82
	mem[16'h463] = 24'h215982; //000034bae
	mem[16'h464] = 24'h215517; //0000349dd
	mem[16'h465] = 24'h215053; //00003480d
	mem[16'h466] = 24'h214592; //000034640
	mem[16'h467] = 24'h214132; //000034474
	mem[16'h468] = 24'h213675; //0000342ab
	mem[16'h469] = 24'h213219; //0000340e3
	mem[16'h486] = 24'h205761; //0000323c1
	mem[16'h487] = 24'h205338; //00003221a
	mem[16'h864] = 24'h115740; //00001c41c
	mem[16'h865] = 24'h115606; //00001c396
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h470] = 24'h212765; //000033f1d
	mem[16'h471] = 24'h212314; //000033d5a
	mem[16'h472] = 24'h211864; //000033b98
	mem[16'h473] = 24'h211416; //0000339d8
	mem[16'h474] = 24'h210970; //00003381a
	mem[16'h475] = 24'h210526; //00003365e
	mem[16'h476] = 24'h210084; //0000334a4
	mem[16'h477] = 24'h209643; //0000332eb
	mem[16'h478] = 24'h209205; //000033135
	mem[16'h479] = 24'h208768; //000032f80
	mem[16'h496] = 24'h201612; //00003138c
	mem[16'h497] = 24'h201207; //0000311f7
	mem[16'h874] = 24'h114416; //00001bef0
	mem[16'h875] = 24'h114285; //00001be6d
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h500] = 24'h200000; //000030d40
	mem[16'h501] = 24'h199600; //000030bb0
	mem[16'h502] = 24'h199203; //000030a23
	mem[16'h503] = 24'h198807; //000030897
	mem[16'h504] = 24'h198412; //00003070c
	mem[16'h505] = 24'h198019; //000030583
	mem[16'h506] = 24'h197628; //0000303fc
	mem[16'h507] = 24'h197238; //000030276
	mem[16'h508] = 24'h196850; //0000300f2
	mem[16'h509] = 24'h196463; //00002ff6f
	mem[16'h580] = 24'h172413; //00002a17d
	mem[16'h581] = 24'h172117; //00002a055
	mem[16'h904] = 24'h110619; //00001b01b
	mem[16'h905] = 24'h110497; //00001afa1
	mem[16'h984] = 24'h101626; //000018cfa
	mem[16'h985] = 24'h101522; //000018c92
	mem[16'h510] = 24'h196078; //00002fdee
	mem[16'h511] = 24'h195694; //00002fc6e
	mem[16'h512] = 24'h195312; //00002faf0
	mem[16'h513] = 24'h194931; //00002f973
	mem[16'h514] = 24'h194552; //00002f7f8
	mem[16'h515] = 24'h194174; //00002f67e
	mem[16'h516] = 24'h193798; //00002f506
	mem[16'h517] = 24'h193423; //00002f38f
	mem[16'h518] = 24'h193050; //00002f21a
	mem[16'h519] = 24'h192678; //00002f0a6
	mem[16'h590] = 24'h169491; //000029613
	mem[16'h591] = 24'h169204; //0000294f4
	mem[16'h914] = 24'h109409; //00001ab61
	mem[16'h915] = 24'h109289; //00001aae9
	mem[16'h994] = 24'h100603; //0000188fb
	mem[16'h995] = 24'h100502; //000018896
	mem[16'h520] = 24'h192307; //00002ef33
	mem[16'h521] = 24'h191938; //00002edc2
	mem[16'h522] = 24'h191570; //00002ec52
	mem[16'h523] = 24'h191204; //00002eae4
	mem[16'h524] = 24'h190839; //00002e977
	mem[16'h525] = 24'h190476; //00002e80c
	mem[16'h526] = 24'h190114; //00002e6a2
	mem[16'h527] = 24'h189753; //00002e539
	mem[16'h528] = 24'h189393; //00002e3d1
	mem[16'h529] = 24'h189035; //00002e26b
	mem[16'h582] = 24'h171821; //000029f2d
	mem[16'h583] = 24'h171526; //000029e06
	mem[16'h924] = 24'h108225; //00001a6c1
	mem[16'h925] = 24'h108108; //00001a64c
	mem[16'h948] = 24'h105485; //000019c0d
	mem[16'h949] = 24'h105374; //000019b9e
	mem[16'h530] = 24'h188679; //00002e107
	mem[16'h531] = 24'h188323; //00002dfa3
	mem[16'h532] = 24'h187969; //00002de41
	mem[16'h533] = 24'h187617; //00002dce1
	mem[16'h534] = 24'h187265; //00002db81
	mem[16'h535] = 24'h186915; //00002da23
	mem[16'h536] = 24'h186567; //00002d8c7
	mem[16'h537] = 24'h186219; //00002d76b
	mem[16'h538] = 24'h185873; //00002d611
	mem[16'h539] = 24'h185528; //00002d4b8
	mem[16'h592] = 24'h168918; //0000293d6
	mem[16'h593] = 24'h168634; //0000292ba
	mem[16'h934] = 24'h107066; //00001a23a
	mem[16'h935] = 24'h106951; //00001a1c7
	mem[16'h958] = 24'h104384; //0000197c0
	mem[16'h959] = 24'h104275; //000019753
	mem[16'h540] = 24'h185185; //00002d361
	mem[16'h541] = 24'h184842; //00002d20a
	mem[16'h542] = 24'h184501; //00002d0b5
	mem[16'h543] = 24'h184162; //00002cf62
	mem[16'h544] = 24'h183823; //00002ce0f
	mem[16'h545] = 24'h183486; //00002ccbe
	mem[16'h546] = 24'h183150; //00002cb6e
	mem[16'h547] = 24'h182815; //00002ca1f
	mem[16'h548] = 24'h182481; //00002c8d1
	mem[16'h549] = 24'h182149; //00002c785
	mem[16'h584] = 24'h171232; //000029ce0
	mem[16'h585] = 24'h170940; //000029bbc
	mem[16'h944] = 24'h105932; //000019dcc
	mem[16'h945] = 24'h105820; //000019d5c
	mem[16'h588] = 24'h170068; //000029854
	mem[16'h589] = 24'h169779; //000029733
	mem[16'h550] = 24'h181818; //00002c63a
	mem[16'h551] = 24'h181488; //00002c4f0
	mem[16'h552] = 24'h181159; //00002c3a7
	mem[16'h553] = 24'h180831; //00002c25f
	mem[16'h554] = 24'h180505; //00002c119
	mem[16'h555] = 24'h180180; //00002bfd4
	mem[16'h556] = 24'h179856; //00002be90
	mem[16'h557] = 24'h179533; //00002bd4d
	mem[16'h558] = 24'h179211; //00002bc0b
	mem[16'h559] = 24'h178890; //00002baca
	mem[16'h594] = 24'h168350; //00002919e
	mem[16'h595] = 24'h168067; //000029083
	mem[16'h954] = 24'h104821; //000019975
	mem[16'h955] = 24'h104712; //000019908
	mem[16'h598] = 24'h167224; //000028d38
	mem[16'h599] = 24'h166944; //000028c20
	mem[16'h560] = 24'h178571; //00002b98b
	mem[16'h561] = 24'h178253; //00002b84d
	mem[16'h562] = 24'h177935; //00002b70f
	mem[16'h563] = 24'h177619; //00002b5d3
	mem[16'h564] = 24'h177304; //00002b498
	mem[16'h565] = 24'h176991; //00002b35f
	mem[16'h566] = 24'h176678; //00002b226
	mem[16'h567] = 24'h176366; //00002b0ee
	mem[16'h568] = 24'h176056; //00002afb8
	mem[16'h569] = 24'h175746; //00002ae82
	mem[16'h586] = 24'h170648; //000029a98
	mem[16'h587] = 24'h170357; //000029975
	mem[16'h964] = 24'h103734; //000019536
	mem[16'h965] = 24'h103626; //0000194ca
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h570] = 24'h175438; //00002ad4e
	mem[16'h571] = 24'h175131; //00002ac1b
	mem[16'h572] = 24'h174825; //00002aae9
	mem[16'h573] = 24'h174520; //00002a9b8
	mem[16'h574] = 24'h174216; //00002a888
	mem[16'h575] = 24'h173913; //00002a759
	mem[16'h576] = 24'h173611; //00002a62b
	mem[16'h577] = 24'h173310; //00002a4fe
	mem[16'h578] = 24'h173010; //00002a3d2
	mem[16'h579] = 24'h172711; //00002a2a7
	mem[16'h596] = 24'h167785; //000028f69
	mem[16'h597] = 24'h167504; //000028e50
	mem[16'h974] = 24'h102669; //00001910d
	mem[16'h975] = 24'h102564; //0000190a4
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h000] = 24'h000000; //000000000
	mem[16'h600] = 24'h166666; //000028b0a
	mem[16'h601] = 24'h166389; //0000289f5
	mem[16'h602] = 24'h166112; //0000288e0
	mem[16'h603] = 24'h165837; //0000287cd
	mem[16'h604] = 24'h165562; //0000286ba
	mem[16'h605] = 24'h165289; //0000285a9
	mem[16'h606] = 24'h165016; //000028498
	mem[16'h607] = 24'h164744; //000028388
	mem[16'h608] = 24'h164473; //000028279
	mem[16'h609] = 24'h164203; //00002816b
	mem[16'h680] = 24'h147058; //000023e72
	mem[16'h681] = 24'h146842; //000023d9a
	mem[16'h806] = 24'h124069; //00001e4a5
	mem[16'h807] = 24'h123915; //00001e40b
	mem[16'h886] = 24'h112866; //00001b8e2
	mem[16'h887] = 24'h112739; //00001b863
	mem[16'h610] = 24'h163934; //00002805e
	mem[16'h611] = 24'h163666; //000027f52
	mem[16'h612] = 24'h163398; //000027e46
	mem[16'h613] = 24'h163132; //000027d3c
	mem[16'h614] = 24'h162866; //000027c32
	mem[16'h615] = 24'h162601; //000027b29
	mem[16'h616] = 24'h162337; //000027a21
	mem[16'h617] = 24'h162074; //00002791a
	mem[16'h618] = 24'h161812; //000027814
	mem[16'h619] = 24'h161550; //00002770e
	mem[16'h690] = 24'h144927; //00002361f
	mem[16'h691] = 24'h144717; //00002354d
	mem[16'h816] = 24'h122549; //00001deb5
	mem[16'h817] = 24'h122399; //00001de1f
	mem[16'h896] = 24'h111607; //00001b3f7
	mem[16'h897] = 24'h111482; //00001b37a
	mem[16'h620] = 24'h161290; //00002760a
	mem[16'h621] = 24'h161030; //000027506
	mem[16'h622] = 24'h160771; //000027403
	mem[16'h623] = 24'h160513; //000027301
	mem[16'h624] = 24'h160256; //000027200
	mem[16'h625] = 24'h160000; //000027100
	mem[16'h626] = 24'h159744; //000027000
	mem[16'h627] = 24'h159489; //000026f01
	mem[16'h628] = 24'h159235; //000026e03
	mem[16'h629] = 24'h158982; //000026d06
	mem[16'h682] = 24'h146627; //000023cc3
	mem[16'h683] = 24'h146412; //000023bec
	mem[16'h826] = 24'h121065; //00001d8e9
	mem[16'h827] = 24'h120918; //00001d856
	mem[16'h868] = 24'h115207; //00001c207
	mem[16'h869] = 24'h115074; //00001c182
	mem[16'h630] = 24'h158730; //000026c0a
	mem[16'h631] = 24'h158478; //000026b0e
	mem[16'h632] = 24'h158227; //000026a13
	mem[16'h633] = 24'h157977; //000026919
	mem[16'h634] = 24'h157728; //000026820
	mem[16'h635] = 24'h157480; //000026728
	mem[16'h636] = 24'h157232; //000026630
	mem[16'h637] = 24'h156985; //000026539
	mem[16'h638] = 24'h156739; //000026443
	mem[16'h639] = 24'h156494; //00002634e
	mem[16'h692] = 24'h144508; //00002347c
	mem[16'h693] = 24'h144300; //0000233ac
	mem[16'h836] = 24'h119617; //00001d341
	mem[16'h837] = 24'h119474; //00001d2b2
	mem[16'h878] = 24'h113895; //00001bce7
	mem[16'h879] = 24'h113765; //00001bc65
	mem[16'h640] = 24'h156250; //00002625a
	mem[16'h641] = 24'h156006; //000026166
	mem[16'h642] = 24'h155763; //000026073
	mem[16'h643] = 24'h155520; //000025f80
	mem[16'h644] = 24'h155279; //000025e8f
	mem[16'h645] = 24'h155038; //000025d9e
	mem[16'h646] = 24'h154798; //000025cae
	mem[16'h647] = 24'h154559; //000025bbf
	mem[16'h648] = 24'h154320; //000025ad0
	mem[16'h649] = 24'h154083; //0000259e3
	mem[16'h684] = 24'h146198; //000023b16
	mem[16'h685] = 24'h145985; //000023a41
	mem[16'h846] = 24'h118203; //00001cdbb
	mem[16'h847] = 24'h118063; //00001cd2f
	mem[16'h688] = 24'h145348; //0000237c4
	mem[16'h689] = 24'h145137; //0000236f1
	mem[16'h650] = 24'h153846; //0000258f6
	mem[16'h651] = 24'h153609; //000025809
	mem[16'h652] = 24'h153374; //00002571e
	mem[16'h653] = 24'h153139; //000025633
	mem[16'h654] = 24'h152905; //000025549
	mem[16'h655] = 24'h152671; //00002545f
	mem[16'h656] = 24'h152439; //000025377
	mem[16'h657] = 24'h152207; //00002528f
	mem[16'h658] = 24'h151975; //0000251a7
	mem[16'h659] = 24'h151745; //0000250c1
	mem[16'h694] = 24'h144092; //0000232dc
	mem[16'h695] = 24'h143884; //00002320c
	mem[16'h856] = 24'h116822; //00001c856
	mem[16'h857] = 24'h116686; //00001c7ce
	mem[16'h698] = 24'h143266; //000022fa2
	mem[16'h699] = 24'h143061; //000022ed5
	mem[16'h660] = 24'h151515; //000024fdb
	mem[16'h661] = 24'h151285; //000024ef5
	mem[16'h662] = 24'h151057; //000024e11
	mem[16'h663] = 24'h150829; //000024d2d
	mem[16'h664] = 24'h150602; //000024c4a
	mem[16'h665] = 24'h150375; //000024b67
	mem[16'h666] = 24'h150150; //000024a86
	mem[16'h667] = 24'h149925; //0000249a5
	mem[16'h668] = 24'h149700; //0000248c4
	mem[16'h669] = 24'h149476; //0000247e4
	mem[16'h686] = 24'h145772; //00002396c
	mem[16'h687] = 24'h145560; //000023898
	mem[16'h866] = 24'h115473; //00001c311
	mem[16'h867] = 24'h115340; //00001c28c
	mem[16'hfff] = 24'hffffff; //fffffffff
	mem[16'hfff] = 24'hffffff; //fffffffff
	mem[16'h670] = 24'h149253; //000024705
	mem[16'h671] = 24'h149031; //000024627
	mem[16'h672] = 24'h148809; //000024549
	mem[16'h673] = 24'h148588; //00002446c
	mem[16'h674] = 24'h148367; //00002438f
	mem[16'h675] = 24'h148148; //0000242b4
	mem[16'h676] = 24'h147928; //0000241d8
	mem[16'h677] = 24'h147710; //0000240fe
	mem[16'h678] = 24'h147492; //000024024
	mem[16'h679] = 24'h147275; //000023f4b
	mem[16'h696] = 24'h143678; //00002313e
	mem[16'h697] = 24'h143472; //000023070
	mem[16'h876] = 24'h114155; //00001bdeb
	mem[16'h877] = 24'h114025; //00001bd69
	mem[16'hfff] = 24'hffffff; //fffffffff
	mem[16'hfff] = 24'hffffff; //fffffffff
	mem[16'h700] = 24'h142857; //000022e09
	mem[16'h701] = 24'h142653; //000022d3d
	mem[16'h702] = 24'h142450; //000022c72
	mem[16'h703] = 24'h142247; //000022ba7
	mem[16'h704] = 24'h142045; //000022add
	mem[16'h705] = 24'h141843; //000022a13
	mem[16'h706] = 24'h141643; //00002294b
	mem[16'h707] = 24'h141442; //000022882
	mem[16'h708] = 24'h141242; //0000227ba
	mem[16'h709] = 24'h141043; //0000226f3
	mem[16'h780] = 24'h128205; //00001f4cd
	mem[16'h781] = 24'h128040; //00001f428
	mem[16'h906] = 24'h110375; //00001af27
	mem[16'h907] = 24'h110253; //00001aead
	mem[16'h986] = 24'h101419; //000018c2b
	mem[16'h987] = 24'h101317; //000018bc5
	mem[16'h710] = 24'h140845; //00002262d
	mem[16'h711] = 24'h140646; //000022566
	mem[16'h712] = 24'h140449; //0000224a1
	mem[16'h713] = 24'h140252; //0000223dc
	mem[16'h714] = 24'h140056; //000022318
	mem[16'h715] = 24'h139860; //000022254
	mem[16'h716] = 24'h139664; //000022190
	mem[16'h717] = 24'h139470; //0000220ce
	mem[16'h718] = 24'h139275; //00002200b
	mem[16'h719] = 24'h139082; //000021f4a
	mem[16'h790] = 24'h126582; //00001ee76
	mem[16'h791] = 24'h126422; //00001edd6
	mem[16'h916] = 24'h109170; //00001aa72
	mem[16'h917] = 24'h109051; //00001a9fb
	mem[16'h996] = 24'h100401; //000018831
	mem[16'h997] = 24'h100300; //0000187cc
	mem[16'h720] = 24'h138888; //000021e88
	mem[16'h721] = 24'h138696; //000021dc8
	mem[16'h722] = 24'h138504; //000021d08
	mem[16'h723] = 24'h138312; //000021c48
	mem[16'h724] = 24'h138121; //000021b89
	mem[16'h725] = 24'h137931; //000021acb
	mem[16'h726] = 24'h137741; //000021a0d
	mem[16'h727] = 24'h137551; //00002194f
	mem[16'h728] = 24'h137362; //000021892
	mem[16'h729] = 24'h137174; //0000217d6
	mem[16'h782] = 24'h127877; //00001f385
	mem[16'h783] = 24'h127713; //00001f2e1
	mem[16'h926] = 24'h107991; //00001a5d7
	mem[16'h927] = 24'h107874; //00001a562
	mem[16'h968] = 24'h103305; //000019389
	mem[16'h969] = 24'h103199; //00001931f
	mem[16'h730] = 24'h136986; //00002171a
	mem[16'h731] = 24'h136798; //00002165e
	mem[16'h732] = 24'h136612; //0000215a4
	mem[16'h733] = 24'h136425; //0000214e9
	mem[16'h734] = 24'h136239; //00002142f
	mem[16'h735] = 24'h136054; //000021376
	mem[16'h736] = 24'h135869; //0000212bd
	mem[16'h737] = 24'h135685; //000021205
	mem[16'h738] = 24'h135501; //00002114d
	mem[16'h739] = 24'h135317; //000021095
	mem[16'h792] = 24'h126262; //00001ed36
	mem[16'h793] = 24'h126103; //00001ec97
	mem[16'h936] = 24'h106837; //00001a155
	mem[16'h937] = 24'h106723; //00001a0e3
	mem[16'h978] = 24'h102249; //000018f69
	mem[16'h979] = 24'h102145; //000018f01
	mem[16'h740] = 24'h135135; //000020fdf
	mem[16'h741] = 24'h134952; //000020f28
	mem[16'h742] = 24'h134770; //000020e72
	mem[16'h743] = 24'h134589; //000020dbd
	mem[16'h744] = 24'h134408; //000020d08
	mem[16'h745] = 24'h134228; //000020c54
	mem[16'h746] = 24'h134048; //000020ba0
	mem[16'h747] = 24'h133868; //000020aec
	mem[16'h748] = 24'h133689; //000020a39
	mem[16'h749] = 24'h133511; //000020987
	mem[16'h784] = 24'h127551; //00001f23f
	mem[16'h785] = 24'h127388; //00001f19c
	mem[16'h946] = 24'h105708; //000019cec
	mem[16'h947] = 24'h105596; //000019c7c
	mem[16'h788] = 24'h126903; //00001efb7
	mem[16'h789] = 24'h126742; //00001ef16
	mem[16'h750] = 24'h133333; //0000208d5
	mem[16'h751] = 24'h133155; //000020823
	mem[16'h752] = 24'h132978; //000020772
	mem[16'h753] = 24'h132802; //0000206c2
	mem[16'h754] = 24'h132625; //000020611
	mem[16'h755] = 24'h132450; //000020562
	mem[16'h756] = 24'h132275; //0000204b3
	mem[16'h757] = 24'h132100; //000020404
	mem[16'h758] = 24'h131926; //000020356
	mem[16'h759] = 24'h131752; //0000202a8
	mem[16'h794] = 24'h125944; //00001ebf8
	mem[16'h795] = 24'h125786; //00001eb5a
	mem[16'h956] = 24'h104602; //00001989a
	mem[16'h957] = 24'h104493; //00001982d
	mem[16'h798] = 24'h125313; //00001e981
	mem[16'h799] = 24'h125156; //00001e8e4
	mem[16'h760] = 24'h131578; //0000201fa
	mem[16'h761] = 24'h131406; //00002014e
	mem[16'h762] = 24'h131233; //0000200a1
	mem[16'h763] = 24'h131061; //00001fff5
	mem[16'h764] = 24'h130890; //00001ff4a
	mem[16'h765] = 24'h130718; //00001fe9e
	mem[16'h766] = 24'h130548; //00001fdf4
	mem[16'h767] = 24'h130378; //00001fd4a
	mem[16'h768] = 24'h130208; //00001fca0
	mem[16'h769] = 24'h130039; //00001fbf7
	mem[16'h786] = 24'h127226; //00001f0fa
	mem[16'h787] = 24'h127064; //00001f058
	mem[16'h966] = 24'h103519; //00001945f
	mem[16'h967] = 24'h103412; //0000193f4
	mem[16'hfff] = 24'hffffff; //fffffffff
	mem[16'hfff] = 24'hffffff; //fffffffff
	mem[16'h770] = 24'h129870; //00001fb4e
	mem[16'h771] = 24'h129701; //00001faa5
	mem[16'h772] = 24'h129533; //00001f9fd
	mem[16'h773] = 24'h129366; //00001f956
	mem[16'h774] = 24'h129198; //00001f8ae
	mem[16'h775] = 24'h129032; //00001f808
	mem[16'h776] = 24'h128865; //00001f761
	mem[16'h777] = 24'h128700; //00001f6bc
	mem[16'h778] = 24'h128534; //00001f616
	mem[16'h779] = 24'h128369; //00001f571
	mem[16'h796] = 24'h125628; //00001eabc
	mem[16'h797] = 24'h125470; //00001ea1e
	mem[16'h976] = 24'h102459; //00001903b
	mem[16'h977] = 24'h102354; //000018fd2
	mem[16'hfff] = 24'hffffff; //fffffffff
	mem[16'hfff] = 24'hffffff; //fffffffff
end

always_ff @(posedge clk)
	ndx <= iu.sig[135:124];
always_ff @(posedge clk)
begin
	ou <= iu;
	ou.exp <= 14'h17FF;
	ou.sig <= {mem[ndx],112'd0};
end

DFPPack128 u2 (ou, o);

endmodule
